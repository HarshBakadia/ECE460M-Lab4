`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: UT Austin
// Engineer: Brandon King
// 
// Create Date: 02/28/2024 05:48:53 PM
// Design Name: Parking Meter
// Module Name: Clk_Gen
// Project Name: Lab 4
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// 1 Pulse of 100MHz every Sec 
module Pulser_1Hz(SYS_CLK, Pulse);
  input SYS_CLK; //fast clock
  output reg Pulse; //slow clock

  reg[27:0] counter;

  initial begin
    counter = 0;
    Pulse = 0;
  end

  always @ (posedge SYS_CLK)
  begin
    if(counter == 100000000) begin
      counter <= 1;
      Pulse <= 'b1;
    end
    else begin
      counter <= counter + 1;
      Pulse <= 'b0;
    end
  end
endmodule

// 1 Pulse/Sec 
module Divider_1Hz(SYS_CLK, slowClk);
  input SYS_CLK; //fast clock
  output reg slowClk; //slow clock

  reg[27:0] counter;

  initial begin
    counter = 0;
    slowClk = 0;
  end

  always @ (posedge SYS_CLK)
  begin
    if(counter == 50000000) begin
      counter <= 1;
      slowClk <= ~slowClk;
    end
    else begin
      counter <= counter + 1;
    end
  end
endmodule


// 15 Pulse/Sec
module Divider_15Hz(SYS_CLK, slowClk);
  input SYS_CLK; //fast clock
  output reg slowClk; //slow clock

  reg[27:0] counter;

  initial begin
    counter = 0;
    slowClk = 0;
  end

  always @ (posedge SYS_CLK)
  begin
    if(counter == 7500000) begin
      counter <= 1;
      slowClk <= ~slowClk;
    end
    else begin
      counter <= counter + 1;
    end
  end
endmodule

// 30kHz Pulse/Sec 
module Divider_30kHz(SYS_CLK, slowClk);
  input SYS_CLK; //fast clock
  output reg slowClk; //slow clock

  reg[27:0] counter;

  initial begin
    counter = 0;
    slowClk = 0;
  end

  always @ (posedge SYS_CLK)
  begin
    if(counter == 00001667) begin
      counter <= 1;
      slowClk <= ~slowClk;
    end
    else begin
      counter <= counter + 1;
    end
  end
endmodule